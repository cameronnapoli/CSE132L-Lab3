module hazardunit(
    output logic StallF,
    output logic StallID,
    output logic FlushID,
    output logic FlushE,
    output logic [1:0] ForwardAE,
    output logic [1:0] ForwardBE,
    output logic Match, // Input or Output ????
    output logic RegWriteM,
    output logic RegWriteW,
    output logic MemtoRegE
    );

endmodule
