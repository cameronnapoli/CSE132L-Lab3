module hazardunit(
    output logic StallF,
    output logic StallID,
    output logic FlushID,
    output logic FlushE,
    output logic ForwardAE,
    output logic ForwardBE,
    output logic Match, // Input or Output ???
    output logic RegWriteM,
    output logic RegWriteW,
    output logic MemtoRegE
    );

endmodule
