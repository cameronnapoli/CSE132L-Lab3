module regIFID(
    input logic clk
    );

endmodule


module regIDEX(
    input logic clk
    );

endmodule


module regEXMEM(
    input logic clk
    );

endmodule


module regMEMWB(
    input logic clk
    );

endmodule
