module mux2
    #(parameter WIDTH = 8)
    (input logic [WIDTH-1:0] d0, d1, d3,
    input logic [1:0] s,
    output logic [WIDTH-1:0] y);

    // Logic for 3 input mux here

endmodule
